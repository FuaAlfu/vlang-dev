module two

// an export  function we have to use `pub` to use it
pub fn hit(a int, b int){
	//I love you)
	println(a-b)
}