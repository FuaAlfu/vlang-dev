module three

// an export  function we have to use `pub` to use it
pub fn three(){
	//I love you)
	println('ya lublu tebya!!')
}