module da

// an export  function we have to use `pub` to use it
pub fn da(){
	//I love you)
	println('ya lublu tebya!!')
}