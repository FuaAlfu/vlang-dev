module one

// an export  function we have to use `pub` to use it
pub fn sum (a int,b int) int{
	
	return a + b
}