module hi

// an export  function we have to use `pub` to use it
pub fn say_hi() {
    println('yo from hi!')
}