const (
	pi    = 3.14
	golden_ratio = 1.6180
)

fn main() {
	/*
	Constants are declared with const keyword.
	They can only be defined at the module level (outside of functions).
	Constant values can never be changed.
	we can also declare a single constant separately
	*/
	println(pi)
    println(golden_ratio)
}

